package imdct_simple_pkg;
  import uvm_pkg::*;      // import the UVM library
  `include "uvm_macros.svh" // Include the UVM macros
  `include "imdct_item.sv"
  `include "imdct_sequencer.sv"

endpackage 