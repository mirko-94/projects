----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 08/24/2022 03:24:06 PM
-- Design Name: 
-- Module Name: cos_rom_1 - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity cos_rom_1 is
    generic (
	       WIDTH : integer := 32;
	       WIDTH_2 : integer := 64;
	       WIDTH_3 : integer := 96; 
	       WADDR   : integer := 8
    );
    port(
        address_cos_1 : in  std_logic_vector(WADDR-1 downto 0);
        dout_cos_1    : out std_logic_vector(WIDTH-1 downto 0)
    );
end cos_rom_1;

architecture Behavioral of cos_rom_1 is
  type mem is array ( 0 to 215) of std_logic_vector(WIDTH-1 downto 0);
  constant my_Rom : mem := (
  
0 => "00111111000110111101011111000011",
1 => "10111111011011001000001101100110",
2 => "10111110000001011010100010011100",
3 => "00111111011111011100111101010111",
4 => "10111110110000111110111100000111",
5 => "10111111010010110001100100101111",
6 => "00111110110000111110111100000111",
7 => "10111111011011001000001101100110",
8 => "00111111011011001000001101100110",
9 => "10111110110000111110111100000111",
10 => "10111110110000111110111100000111",
11 => "00111111011011001000001101100110",
12 => "00111110000001011010100010011100",
13 => "10111110110000111110111100000111",
14 => "00111111000110111101011111000011",
15 => "10111111010010110001100100101111",
16 => "00111111011011001000001101100110",
17 => "10111111011111011100111101010111",
18 => "10111110000001011010100010011100",
19 => "00111110110000111110111100000111",
20 => "10111111000110111101011111000011",
21 => "00111111010010110001100100101111",
22 => "10111111011011001000001101100110",
23 => "00111111011111011100111101010111",
24 => "10111110110000111110111100000111",
25 => "00111111011011001000001101100110",
26 => "10111111011011001000001101100110",
27 => "00111110110000111110111100000111",
28 => "00111110110000111110111100000111",
29 => "10111111011011001000001101100110",
30 => "10111111000110111101011111000011",
31 => "00111111011011001000001101100110",
32 => "00111110000001011010100010011100",
33 => "10111111011111011100111101010111",
34 => "00111110110000111110111100000111",
35 => "00111111010010110001100100101111",
36 => "10111111010010110001100100101111",
37 => "00111110110000111110111100000111",
38 => "00111111011111011100111101010111",
39 => "00111110000001011010100010011100",
40 => "10111111011011001000001101100110",
41 => "10111111000110111101011111000011",
42 => "10111111011011001000001101100110",
43 => "10111110110000111110111100000111",
44 => "00111110110000111110111100000111",
45 => "00111111011011001000001101100110",
46 => "00111111011011001000001101100110",
47 => "00111110110000111110111100000111",
48 => "10111111011111011100111101010111",
49 => "10111111011011001000001101100110",
50 => "10111111010010110001100100101111",
51 => "10111111000110111101011111000011",
52 => "10111110110000111110111100000111",
53 => "10111110000001011010100010011100",
54 => "10111111011111011100111101010111",
55 => "10111111011011001000001101100110",
56 => "10111111010010110001100100101111",
57 => "10111111000110111101011111000011",
58 => "10111110110000111110111100000111",
59 => "10111110000001011010100010011100",
60 => "10111111011011001000001101100110",
61 => "10111110110000111110111100000111",
62 => "00111110110000111110111100000111",
63 => "00111111011011001000001101100110",
64 => "00111111011011001000001101100110",
65 => "00111110110000111110111100000111",
66 => "10111111010010110001100100101111",
67 => "00111110110000111110111100000111",
68 => "00111111011111011100111101010111",
69 => "00111110000001011010100010011100",
70 => "10111111011011001000001101100110",
71 => "10111111000110111101011111000011",
72 => "00111111000110111101011111000011",
73 => "10111111011011001000001101100110",
74 => "10111110000001011010100010011100",
75 => "00111111011111011100111101010111",
76 => "10111110110000111110111100000111",
77 => "10111111010010110001100100101111",
78 => "00111110110000111110111100000111",
79 => "10111111011011001000001101100110",
80 => "00111111011011001000001101100110",
81 => "10111110110000111110111100000111",
82 => "10111110110000111110111100000111",
83 => "00111111011011001000001101100110",
84 => "00111110000001011010100010011100",
85 => "10111110110000111110111100000111",
86 => "00111111000110111101011111000011",
87 => "10111111010010110001100100101111",
88 => "00111111011011001000001101100110",
89 => "10111111011111011100111101010111",
90 => "10111110000001011010100010011100",
91 => "00111110110000111110111100000111",
92 => "10111111000110111101011111000011",
93 => "00111111010010110001100100101111",
94 => "10111111011011001000001101100110",
95 => "00111111011111011100111101010111",
96 => "10111110110000111110111100000111",
97 => "00111111011011001000001101100110",
98 => "10111111011011001000001101100110",
99 => "00111110110000111110111100000111",
100 => "00111110110000111110111100000111",
101 => "10111111011011001000001101100110",
102 => "10111111000110111101011111000011",
103 => "00111111011011001000001101100110",
104 => "00111110000001011010100010011100",
105 => "10111111011111011100111101010111",
106 => "00111110110000111110111100000111",
107 => "00111111010010110001100100101111",
108 => "10111111010010110001100100101111",
109 => "00111110110000111110111100000111",
110 => "00111111011111011100111101010111",
111 => "00111110000001011010100010011100",
112 => "10111111011011001000001101100110",
113 => "10111111000110111101011111000011",
114 => "10111111011011001000001101100110",
115 => "10111110110000111110111100000111",
116 => "00111110110000111110111100000111",
117 => "00111111011011001000001101100110",
118 => "00111111011011001000001101100110",
119 => "00111110110000111110111100000111",
120 => "10111111011111011100111101010111",
121 => "10111111011011001000001101100110",
122 => "10111111010010110001100100101111",
123 => "10111111000110111101011111000011",
124 => "10111110110000111110111100000111",
125 => "10111110000001011010100010011100",
126 => "10111111011111011100111101010111",
127 => "10111111011011001000001101100110",
128 => "10111111010010110001100100101111",
129 => "10111111000110111101011111000011",
130 => "10111110110000111110111100000111",
131 => "10111110000001011010100010011100",
132 => "10111111011011001000001101100110",
133 => "10111110110000111110111100000111",
134 => "00111110110000111110111100000111",
135 => "00111111011011001000001101100110",
136 => "00111111011011001000001101100110",
137 => "00111110110000111110111100000111",
138 => "10111111010010110001100100101111",
139 => "00111110110000111110111100000111",
140 => "00111111011111011100111101010111",
141 => "00111110000001011010100010011100",
142 => "10111111011011001000001101100110",
143 => "10111111000110111101011111000011",
144 => "00111111000110111101011111000011",
145 => "10111111011011001000001101100110",
146 => "10111110000001011010100010011100",
147 => "00111111011111011100111101010111",
148 => "10111110110000111110111100000111",
149 => "10111111010010110001100100101111",
150 => "00111110110000111110111100000111",
151 => "10111111011011001000001101100110",
152 => "00111111011011001000001101100110",
153 => "10111110110000111110111100000111",
154 => "10111110110000111110111100000111",
155 => "00111111011011001000001101100110",
156 => "00111110000001011010100010011100",
157 => "10111110110000111110111100000111",
158 => "00111111000110111101011111000011",
159 => "10111111010010110001100100101111",
160 => "00111111011011001000001101100110",
161 => "10111111011111011100111101010111",
162 => "10111110000001011010100010011100",
163 => "00111110110000111110111100000111",
164 => "10111111000110111101011111000011",
165 => "00111111010010110001100100101111",
166 => "10111111011011001000001101100110",
167 => "00111111011111011100111101010111",
168 => "10111110110000111110111100000111",
169 => "00111111011011001000001101100110",
170 => "10111111011011001000001101100110",
171 => "00111110110000111110111100000111",
172 => "00111110110000111110111100000111",
173 => "10111111011011001000001101100110",
174 => "10111111000110111101011111000011",
175 => "00111111011011001000001101100110",
176 => "00111110000001011010100010011100",
177 => "10111111011111011100111101010111",
178 => "00111110110000111110111100000111",
179 => "00111111010010110001100100101111",
180 => "10111111010010110001100100101111",
181 => "00111110110000111110111100000111",
182 => "00111111011111011100111101010111",
183 => "00111110000001011010100010011100",
184 => "10111111011011001000001101100110",
185 => "10111111000110111101011111000011",
186 => "10111111011011001000001101100110",
187 => "10111110110000111110111100000111",
188 => "00111110110000111110111100000111",
189 => "00111111011011001000001101100110",
190 => "00111111011011001000001101100110",
191 => "00111110110000111110111100000111",
192 => "10111111011111011100111101010111",
193 => "10111111011011001000001101100110",
194 => "10111111010010110001100100101111",
195 => "10111111000110111101011111000011",
196 => "10111110110000111110111100000111",
197 => "10111110000001011010100010011100",
198 => "10111111011111011100111101010111",
199 => "10111111011011001000001101100110",
200 => "10111111010010110001100100101111",
201 => "10111111000110111101011111000011",
202 => "10111110110000111110111100000111",
203 => "10111110000001011010100010011100",
204 => "10111111011011001000001101100110",
205 => "10111110110000111110111100000111",
206 => "00111110110000111110111100000111",
207 => "00111111011011001000001101100110",
208 => "00111111011011001000001101100110",
209 => "00111110110000111110111100000111",
210 => "10111111010010110001100100101111",
211 => "00111110110000111110111100000111",
212 => "00111111011111011100111101010111",
213 => "00111110000001011010100010011100",
214 => "10111111011011001000001101100110",
215 => "10111111000110111101011111000011" );
begin

    main : process(address_cos_1)
    begin
        dout_cos_1 <= my_Rom(to_integer(unsigned(address_cos_1)));
    end process main;

end Behavioral;

